`timescale 1ns/1ns
`include "mux16x1.v"

module testbench();
reg [15:0] w;
reg [3:0] s;
wire out;

mux16x1 m(w,s,out);
initial
begin
    $dumpfile("mux16x1.vcd");
    $dumpvars(0,testbench);

    w = 16'b1110100101100101; s=4'b0000;
    #20;

    w = 16'b1110100101100101; s=4'b0001;
    #20;

    w = 16'b1110100101100101; s=4'b0010;
    #20;

    w = 16'b1110100101100101; s=4'b0011;
    #20;

    w = 16'b1110100101100101; s=4'b0100;
    #20;

    w = 16'b1110100101100101; s=4'b0101;
    #20;

    w = 16'b1110100101100101; s=4'b0110;
    #20;

    w = 16'b1110100101100101; s=4'b0111;
    #20;
    
    w = 16'b1110100101100101; s=4'b1000;
    #20;

    w = 16'b1110100101100101; s=4'b1001;
    #20;

    w = 16'b1110100101100101; s=4'b1010;
    #20;

    w = 16'b1110100101100101; s=4'b1011;
    #20;
    
    w = 16'b1110100101100101; s=4'b1100;
    #20;

    w = 16'b1110100101100101; s=4'b1101;
    #20;

    w = 16'b1110100101100101; s=4'b1110;
    #20;

    w = 16'b1110100101100101; s=4'b1111;
    #20;
    
    $display("test complete");
end
endmodule